module lut_u_module #(
    parameter DATA_WIDTH=16,
    parameter ADDR_WIDTH=8
    )(
        input enable,
        input [(ADDR_WIDTH-1):0] addr,
        output reg [(DATA_WIDTH-1):0] q
        );


    always @ ( * ) begin
        if(enable) begin
            case(addr)
                8'd0 : q = 16'd4;
                8'd16 : q = 16'd8;
                8'd17 : q = 16'd4;
                8'd32 : q = 16'd12;
                8'd33 : q = 16'd8;
                8'd34 : q = 16'd4;
                8'd48 : q = 16'd16;
                8'd49 : q = 16'd12;
                8'd50 : q = 16'd8;
                8'd51 : q = 16'd4;
                8'd64 : q = 16'd20;
                8'd65 : q = 16'd16;
                8'd66 : q = 16'd12;
                8'd67 : q = 16'd8;
                8'd68 : q = 16'd4;
                8'd80 : q = 16'd24;
                8'd81 : q = 16'd20;
                8'd82 : q = 16'd16;
                8'd83 : q = 16'd12;
                8'd84 : q = 16'd8;
                8'd85 : q = 16'd4;
                8'd96 : q = 16'd28;
                8'd97 : q = 16'd24;
                8'd98 : q = 16'd20;
                8'd99 : q = 16'd16;
                8'd100 : q = 16'd12;
                8'd101 : q = 16'd8;
                8'd102 : q = 16'd4;
                8'd112 : q = 16'd32;
                8'd113 : q = 16'd28;
                8'd114 : q = 16'd24;
                8'd115 : q = 16'd20;
                8'd116 : q = 16'd16;
                8'd117 : q = 16'd12;
                8'd118 : q = 16'd8;
                8'd119 : q = 16'd4;
                8'd128 : q = 16'd36;
                8'd129 : q = 16'd32;
                8'd130 : q = 16'd28;
                8'd131 : q = 16'd24;
                8'd132 : q = 16'd20;
                8'd133 : q = 16'd16;
                8'd134 : q = 16'd12;
                8'd135 : q = 16'd8;
                8'd136 : q = 16'd4;
                8'd144 : q = 16'd40;
                8'd145 : q = 16'd36;
                8'd146 : q = 16'd32;
                8'd147 : q = 16'd28;
                8'd148 : q = 16'd24;
                8'd149 : q = 16'd20;
                8'd150 : q = 16'd16;
                8'd151 : q = 16'd12;
                8'd152 : q = 16'd8;
                8'd153 : q = 16'd4;
                8'd160 : q = 16'd44;
                8'd161 : q = 16'd40;
                8'd162 : q = 16'd36;
                8'd163 : q = 16'd32;
                8'd164 : q = 16'd28;
                8'd165 : q = 16'd24;
                8'd166 : q = 16'd20;
                8'd167 : q = 16'd16;
                8'd168 : q = 16'd12;
                8'd169 : q = 16'd8;
                8'd170 : q = 16'd4;
                8'd176 : q = 16'd48;
                8'd177 : q = 16'd44;
                8'd178 : q = 16'd40;
                8'd179 : q = 16'd36;
                8'd180 : q = 16'd32;
                8'd181 : q = 16'd28;
                8'd182 : q = 16'd24;
                8'd183 : q = 16'd20;
                8'd184 : q = 16'd16;
                8'd185 : q = 16'd12;
                8'd186 : q = 16'd8;
                8'd187 : q = 16'd4;
                8'd192 : q = 16'd52;
                8'd193 : q = 16'd48;
                8'd194 : q = 16'd44;
                8'd195 : q = 16'd40;
                8'd196 : q = 16'd36;
                8'd197 : q = 16'd32;
                8'd198 : q = 16'd28;
                8'd199 : q = 16'd24;
                8'd200 : q = 16'd20;
                8'd201 : q = 16'd16;
                8'd202 : q = 16'd12;
                8'd203 : q = 16'd8;
                8'd204 : q = 16'd4;
                8'd208 : q = 16'd56;
                8'd209 : q = 16'd52;
                8'd210 : q = 16'd48;
                8'd211 : q = 16'd44;
                8'd212 : q = 16'd40;
                8'd213 : q = 16'd36;
                8'd214 : q = 16'd32;
                8'd215 : q = 16'd28;
                8'd216 : q = 16'd24;
                8'd217 : q = 16'd20;
                8'd218 : q = 16'd16;
                8'd219 : q = 16'd12;
                8'd220 : q = 16'd8;
                8'd221 : q = 16'd4;
                8'd224 : q = 16'd60;
                8'd225 : q = 16'd56;
                8'd226 : q = 16'd52;
                8'd227 : q = 16'd48;
                8'd228 : q = 16'd44;
                8'd229 : q = 16'd40;
                8'd230 : q = 16'd36;
                8'd231 : q = 16'd32;
                8'd232 : q = 16'd28;
                8'd233 : q = 16'd24;
                8'd234 : q = 16'd20;
                8'd235 : q = 16'd16;
                8'd236 : q = 16'd12;
                8'd237 : q = 16'd8;
                8'd238 : q = 16'd4;
                8'd240 : q = 16'd64;
                8'd241 : q = 16'd60;
                8'd242 : q = 16'd56;
                8'd243 : q = 16'd52;
                8'd244 : q = 16'd48;
                8'd245 : q = 16'd44;
                8'd246 : q = 16'd40;
                8'd247 : q = 16'd36;
                8'd248 : q = 16'd32;
                8'd249 : q = 16'd28;
                8'd250 : q = 16'd24;
                8'd251 : q = 16'd20;
                8'd252 : q = 16'd16;
                8'd253 : q = 16'd12;
                8'd254 : q = 16'd8;
                8'd255 : q = 16'd4;
                default: q = 16'd0;
            endcase
        end
    end
endmodule


module lut_v_module #(
    parameter DATA_WIDTH=16,
    parameter ADDR_WIDTH=8
    )(
          input [(ADDR_WIDTH-1):0] addr,
          output reg [(DATA_WIDTH-1):0] q
);

    always @ ( * ) begin
        case(addr)
            8'd16 : q = 16'd4;
            8'd32 : q = 16'd8;
            8'd33 : q = 16'd4;
            8'd48 : q = 16'd12;
            8'd49 : q = 16'd8;
            8'd50 : q = 16'd4;
            8'd64 : q = 16'd16;
            8'd65 : q = 16'd12;
            8'd66 : q = 16'd8;
            8'd67 : q = 16'd4;
            8'd80 : q = 16'd20;
            8'd81 : q = 16'd16;
            8'd82 : q = 16'd12;
            8'd83 : q = 16'd8;
            8'd84 : q = 16'd4;
            8'd96 : q = 16'd24;
            8'd97 : q = 16'd20;
            8'd98 : q = 16'd16;
            8'd99 : q = 16'd12;
            8'd100 : q = 16'd8;
            8'd101 : q = 16'd4;
            8'd112 : q = 16'd28;
            8'd113 : q = 16'd24;
            8'd114 : q = 16'd20;
            8'd115 : q = 16'd16;
            8'd116 : q = 16'd12;
            8'd117 : q = 16'd8;
            8'd118 : q = 16'd4;
            8'd128 : q = 16'd32;
            8'd129 : q = 16'd28;
            8'd130 : q = 16'd24;
            8'd131 : q = 16'd20;
            8'd132 : q = 16'd16;
            8'd133 : q = 16'd12;
            8'd134 : q = 16'd8;
            8'd135 : q = 16'd4;
            8'd144 : q = 16'd36;
            8'd145 : q = 16'd32;
            8'd146 : q = 16'd28;
            8'd147 : q = 16'd24;
            8'd148 : q = 16'd20;
            8'd149 : q = 16'd16;
            8'd150 : q = 16'd12;
            8'd151 : q = 16'd8;
            8'd152 : q = 16'd4;
            8'd160 : q = 16'd40;
            8'd161 : q = 16'd36;
            8'd162 : q = 16'd32;
            8'd163 : q = 16'd28;
            8'd164 : q = 16'd24;
            8'd165 : q = 16'd20;
            8'd166 : q = 16'd16;
            8'd167 : q = 16'd12;
            8'd168 : q = 16'd8;
            8'd169 : q = 16'd4;
            8'd176 : q = 16'd44;
            8'd177 : q = 16'd40;
            8'd178 : q = 16'd36;
            8'd179 : q = 16'd32;
            8'd180 : q = 16'd28;
            8'd181 : q = 16'd24;
            8'd182 : q = 16'd20;
            8'd183 : q = 16'd16;
            8'd184 : q = 16'd12;
            8'd185 : q = 16'd8;
            8'd186 : q = 16'd4;
            8'd192 : q = 16'd48;
            8'd193 : q = 16'd44;
            8'd194 : q = 16'd40;
            8'd195 : q = 16'd36;
            8'd196 : q = 16'd32;
            8'd197 : q = 16'd28;
            8'd198 : q = 16'd24;
            8'd199 : q = 16'd20;
            8'd200 : q = 16'd16;
            8'd201 : q = 16'd12;
            8'd202 : q = 16'd8;
            8'd203 : q = 16'd4;
            8'd208 : q = 16'd52;
            8'd209 : q = 16'd48;
            8'd210 : q = 16'd44;
            8'd211 : q = 16'd40;
            8'd212 : q = 16'd36;
            8'd213 : q = 16'd32;
            8'd214 : q = 16'd28;
            8'd215 : q = 16'd24;
            8'd216 : q = 16'd20;
            8'd217 : q = 16'd16;
            8'd218 : q = 16'd12;
            8'd219 : q = 16'd8;
            8'd220 : q = 16'd4;
            8'd224 : q = 16'd56;
            8'd225 : q = 16'd52;
            8'd226 : q = 16'd48;
            8'd227 : q = 16'd44;
            8'd228 : q = 16'd40;
            8'd229 : q = 16'd36;
            8'd230 : q = 16'd32;
            8'd231 : q = 16'd28;
            8'd232 : q = 16'd24;
            8'd233 : q = 16'd20;
            8'd234 : q = 16'd16;
            8'd235 : q = 16'd12;
            8'd236 : q = 16'd8;
            8'd237 : q = 16'd4;
            8'd240 : q = 16'd60;
            8'd241 : q = 16'd56;
            8'd242 : q = 16'd52;
            8'd243 : q = 16'd48;
            8'd244 : q = 16'd44;
            8'd245 : q = 16'd40;
            8'd246 : q = 16'd36;
            8'd247 : q = 16'd32;
            8'd248 : q = 16'd28;
            8'd249 : q = 16'd24;
            8'd250 : q = 16'd20;
            8'd251 : q = 16'd16;
            8'd252 : q = 16'd12;
            8'd253 : q = 16'd8;
            8'd254 : q = 16'd4;
            default : q = 16'd0;
        endcase
    end
endmodule
