`include "uvm_macros.svh"

`include "header.svh"
`include "top_uvm.sv"
`include "sequence.sv"
`include "driver.sv"
`include "model.sv"
`include "scoreboard.sv"

