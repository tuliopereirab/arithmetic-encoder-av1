`include "uvm_macros.svh"

`include "header.svh"
`include "top_uvm.sv"

//  Module: top_tb
//
module top_tb;
  import uvm_pkg::*;
  import av1_ee_rand_1_bool_uvm::*;
  // TODO
  // 1. interface declaration
  // 2. top_entity declaration & interface connection
  // 3. clk generation
  // 4. Uvm instantiation  
endmodule: top_tb

