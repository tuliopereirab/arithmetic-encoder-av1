module arithmetic_encoder #(
    parameter GENERAL_DATA_16 = 16,
    parameter GENERAL_DATA_32 = 32,
    parameter GENERAL_SYMBOL_WIDTH = 4,
    parameter GENERAL_LUT_ADDR_WIDTH = 8,
    parameter GENERAL_LUT_DATA_WIDTH = 16,
    parameter GENERAL_D_SIZE = 4
    )(
        input general_clk, reset,
        input [(GENERAL_DATA_16-1):0] general_fl, general_fh,
        input [(GENERAL_SYMBOL_WIDTH-1):0] general_symbol,
        input [GENERAL_SYMBOL_WIDTH:0] general_nsyms,
        output wire [(GENERAL_DATA_16-1):0] RANGE_OUTPUT, LOW_OUTPUT,
        output wire [(GENERAL_DATA_32-1):0] CNT_OUTPUT
    );

    // general
    reg [(GENERAL_DATA_16-1):0] reg_Range_s3, reg_Low_s3;
    reg [(GENERAL_DATA_32-1):0] reg_Cnt_s3;
    assign RANGE_OUTPUT = reg_Range_s3;
    assign LOW_OUTPUT = reg_Low_s3;
    assign CNT_OUTPUT = reg_Cnt_s3;

    // control unit
    wire ctrl_reg_1_2, ctrl_reg_2_3, ctrl_reg_final;

    control_unit control (
        .clk (general_clk),
        .reset_ctrl (reset),
        //outputs
        .pipeline_reg_1_2 (ctrl_reg_1_2),
        .pipeline_reg_2_3 (ctrl_reg_2_3),
        .pipeline_reg_final (ctrl_reg_final)
        );


    // stage 1
    wire [(GENERAL_LUT_DATA_WIDTH-1):0] lut_u_output, lut_v_output;
    wire [(GENERAL_DATA_16-1):0] uu_out, vv_out;
    wire COMP_mux_1_out;
    reg [(GENERAL_LUT_DATA_WIDTH-1):0] reg_lut_u, reg_lut_v;
    reg [(GENERAL_DATA_16-1):0] reg_UU, reg_VV;
    reg reg_COMP_mux_1;
    // stage 2
    wire [(GENERAL_DATA_16-1):0] range_out_s2, low_out_s2, mux_reset_range, mux_reset_low;
    reg [(GENERAL_DATA_16-1):0] reg_Range_s2, reg_Low_s2;
    // stage 3, 4, 5
    wire [(GENERAL_DATA_16-1):0] range_out_s3, low_out_s3;
    wire [(GENERAL_DATA_32-1):0] cnt_out_s3;

    // ---------------------------------------------------
    wire [(GENERAL_DATA_16-1):0] init_range, init_low;
    wire [(GENERAL_DATA_32-1):0] init_cnt;
    assign init_range = 16'b1000_0000_0000_0000;                // 16'd32768;
    assign init_low = 16'b0000_0000_0000_0000;                  // 16'd0;
    assign init_cnt = 32'b11111111_11111111_11111111_11110111;  // 32'd4294967287;
    // reset
    always @ (posedge general_clk) begin
        if(reset) begin
            reg_Range_s3 <= init_range;
            reg_Low_s3 <= init_low;
            reg_Cnt_s3 <= init_cnt;
        end
        else if(ctrl_reg_final) begin  // already saving what comes from the Stage [3,4,5]
            reg_Range_s3 <= range_out_s3;
            reg_Low_s3 <= low_out_s3;
            reg_Cnt_s3 <= cnt_out_s3;
        end
    end
    // ---------------------------------------------------
    stage_1 #(
        .DATA_16 (GENERAL_DATA_16),
        .SYMBOL_WIDTH (GENERAL_SYMBOL_WIDTH),
        .LUT_ADDR_WIDTH (GENERAL_LUT_ADDR_WIDTH),
        .LUT_DATA_WIDTH (GENERAL_LUT_DATA_WIDTH)
        ) state_pipeline_1 (
            .clk_stage_1 (general_clk),
            .FL (general_fl),
            .FH (general_fh),
            .SYMBOL (general_symbol),
            .NSYMS (general_nsyms),
            // outputs
            .lut_u_out (lut_u_output),
            .lut_v_out (lut_v_output),
            .UU (uu_out),
            .VV (vv_out),
            .COMP_mux_1 (COMP_mux_1_out)
        );

    always @ (posedge general_clk) begin
        if(ctrl_reg_1_2) begin
            reg_lut_u <= lut_u_output;
            reg_lut_v <= lut_v_output;
            reg_UU <= uu_out;
            reg_VV <= vv_out;
            reg_COMP_mux_1 <= COMP_mux_1_out;
        end
    end
    // ---------------------------------------------------
    stage_2 #(
        .DATA_16 (GENERAL_DATA_16),
        .DATA_32 (GENERAL_DATA_32)
        ) state_pipeline_2 (
            .lut_u (reg_lut_u),
            .lut_v (reg_lut_v),
            .UU (reg_UU),
            .VV (reg_VV),
            .in_range (RANGE_OUTPUT),
            .in_low (LOW_OUTPUT),
            .COMP_mux_1 (reg_COMP_mux_1),
            // outputs
            .range (range_out_s2),
            .low (low_out_s2)
        );

    always @ (posedge general_clk) begin
        if(ctrl_reg_2_3) begin
            reg_Range_s2 <= range_out_s2;
            reg_Low_s2 <= low_out_s2;
        end
    end
    // ---------------------------------------------------
    stage_3_4_5 #(
        .DATA_16 (GENERAL_DATA_16),
        .DATA_32 (GENERAL_DATA_32),
        .D_SIZE (GENERAL_D_SIZE)
        ) state_pipeline_3 (
            .low (reg_Low_s2),
            .range (reg_Range_s2),
            .in_cnt (reg_Cnt_s3),
            // outputs
            .out_low (low_out_s3),
            .out_range (range_out_s3),
            .out_cnt (cnt_out_s3)
        );
endmodule
