module lut_u_module #(
    parameter DATA_WIDTH=16,
    parameter ADDR_WIDTH=8
    )(
          input [(ADDR_WIDTH-1):0] addr,
          output wire [(DATA_WIDTH-1):0] q
);


	assign q = (addr == 0) ? 16'd4 :
               (addr == 16) ? 16'd8 :
               (addr == 17) ? 16'd4 :
               (addr == 32) ? 16'd12 :
               (addr == 33) ? 16'd8 :
               (addr == 34) ? 16'd4 :
               (addr == 48) ? 16'd16 :
               (addr == 49) ? 16'd12 :
               (addr == 50) ? 16'd8 :
               (addr == 51) ? 16'd4 :
               (addr == 64) ? 16'd20 :
               (addr == 65) ? 16'd16 :
               (addr == 66) ? 16'd12 :
               (addr == 67) ? 16'd8 :
               (addr == 68) ? 16'd4 :
               (addr == 80) ? 16'd24 :
               (addr == 81) ? 16'd20 :
               (addr == 82) ? 16'd16 :
               (addr == 83) ? 16'd12 :
               (addr == 84) ? 16'd8 :
               (addr == 85) ? 16'd4 :
               (addr == 96) ? 16'd28 :
               (addr == 97) ? 16'd24 :
               (addr == 98) ? 16'd20 :
               (addr == 99) ? 16'd16 :
               (addr == 100) ? 16'd12 :
               (addr == 101) ? 16'd8 :
               (addr == 102) ? 16'd4 :
               (addr == 112) ? 16'd32 :
               (addr == 113) ? 16'd28 :
               (addr == 114) ? 16'd24 :
               (addr == 115) ? 16'd20 :
               (addr == 116) ? 16'd16 :
               (addr == 117) ? 16'd12 :
               (addr == 118) ? 16'd8 :
               (addr == 119) ? 16'd4 :
               (addr == 128) ? 16'd36 :
               (addr == 129) ? 16'd32 :
               (addr == 130) ? 16'd28 :
               (addr == 131) ? 16'd24 :
               (addr == 132) ? 16'd20 :
               (addr == 133) ? 16'd16 :
               (addr == 134) ? 16'd12 :
               (addr == 135) ? 16'd8 :
               (addr == 136) ? 16'd4 :
               (addr == 144) ? 16'd40 :
               (addr == 145) ? 16'd36 :
               (addr == 146) ? 16'd32 :
               (addr == 147) ? 16'd28 :
               (addr == 148) ? 16'd24 :
               (addr == 149) ? 16'd20 :
               (addr == 150) ? 16'd16 :
               (addr == 151) ? 16'd12 :
               (addr == 152) ? 16'd8 :
               (addr == 153) ? 16'd4 :
               (addr == 160) ? 16'd44 :
               (addr == 161) ? 16'd40 :
               (addr == 162) ? 16'd36 :
               (addr == 163) ? 16'd32 :
               (addr == 164) ? 16'd28 :
               (addr == 165) ? 16'd24 :
               (addr == 166) ? 16'd20 :
               (addr == 167) ? 16'd16 :
               (addr == 168) ? 16'd12 :
               (addr == 169) ? 16'd8 :
               (addr == 170) ? 16'd4 :
               (addr == 176) ? 16'd48 :
               (addr == 177) ? 16'd44 :
               (addr == 178) ? 16'd40 :
               (addr == 179) ? 16'd36 :
               (addr == 180) ? 16'd32 :
               (addr == 181) ? 16'd28 :
               (addr == 182) ? 16'd24 :
               (addr == 183) ? 16'd20 :
               (addr == 184) ? 16'd16 :
               (addr == 185) ? 16'd12 :
               (addr == 186) ? 16'd8 :
               (addr == 187) ? 16'd4 :
               (addr == 192) ? 16'd52 :
               (addr == 193) ? 16'd48 :
               (addr == 194) ? 16'd44 :
               (addr == 195) ? 16'd40 :
               (addr == 196) ? 16'd36 :
               (addr == 197) ? 16'd32 :
               (addr == 198) ? 16'd28 :
               (addr == 199) ? 16'd24 :
               (addr == 200) ? 16'd20 :
               (addr == 201) ? 16'd16 :
               (addr == 202) ? 16'd12 :
               (addr == 203) ? 16'd8 :
               (addr == 204) ? 16'd4 :
               (addr == 208) ? 16'd56 :
               (addr == 209) ? 16'd52 :
               (addr == 210) ? 16'd48 :
               (addr == 211) ? 16'd44 :
               (addr == 212) ? 16'd40 :
               (addr == 213) ? 16'd36 :
               (addr == 214) ? 16'd32 :
               (addr == 215) ? 16'd28 :
               (addr == 216) ? 16'd24 :
               (addr == 217) ? 16'd20 :
               (addr == 218) ? 16'd16 :
               (addr == 219) ? 16'd12 :
               (addr == 220) ? 16'd8 :
               (addr == 221) ? 16'd4 :
               (addr == 224) ? 16'd60 :
               (addr == 225) ? 16'd56 :
               (addr == 226) ? 16'd52 :
               (addr == 227) ? 16'd48 :
               (addr == 228) ? 16'd44 :
               (addr == 229) ? 16'd40 :
               (addr == 230) ? 16'd36 :
               (addr == 231) ? 16'd32 :
               (addr == 232) ? 16'd28 :
               (addr == 233) ? 16'd24 :
               (addr == 234) ? 16'd20 :
               (addr == 235) ? 16'd16 :
               (addr == 236) ? 16'd12 :
               (addr == 237) ? 16'd8 :
               (addr == 238) ? 16'd4 :
               (addr == 240) ? 16'd64 :
               (addr == 241) ? 16'd60 :
               (addr == 242) ? 16'd56 :
               (addr == 243) ? 16'd52 :
               (addr == 244) ? 16'd48 :
               (addr == 245) ? 16'd44 :
               (addr == 246) ? 16'd40 :
               (addr == 247) ? 16'd36 :
               (addr == 248) ? 16'd32 :
               (addr == 249) ? 16'd28 :
               (addr == 250) ? 16'd24 :
               (addr == 251) ? 16'd20 :
               (addr == 252) ? 16'd16 :
               (addr == 253) ? 16'd12 :
               (addr == 254) ? 16'd8 :
               (addr == 255) ? 16'd4 :
               16'd0;


endmodule
