// To check later
// 1- Make the bitstream generation (out_bit_1/2) to be 9-bit arrays

module stage_3 #(
  parameter RANGE_WIDTH = 16,
  parameter LOW_WIDTH = 24,
  parameter D_SIZE = 5
  ) (
    input [(RANGE_WIDTH-1):0] in_range, range_ready, pre_low,
    input [(D_SIZE-1):0] d,
    input COMP_mux_1, bool_flag, symbol,
    input [RANGE_WIDTH:0] u,
    input [(D_SIZE-1):0] in_s,
    input [(LOW_WIDTH-1):0] in_low,
    output wire [(LOW_WIDTH-1):0] out_low,
    output wire [(RANGE_WIDTH-1):0] out_range,
    output wire [(RANGE_WIDTH-1):0] out_bit_1, out_bit_2,
    output wire [1:0] flag_bitstream,
    output wire [(D_SIZE-1):0] out_s
  );
  wire [(LOW_WIDTH-1):0] low_bool, low_cdf;
  wire [(LOW_WIDTH-1):0] low_raw;
  wire [(D_SIZE-1):0] s_bool, s_cdf;
  wire [(RANGE_WIDTH-1):0] out_bit_1_cdf, out_bit_2_cdf;
  wire [(RANGE_WIDTH-1):0] bool_out_bit_1, bool_out_bit_2;
  wire [1:0] flag_cdf, flag_bit_bool;

  s3_cdf #(
    .D_SIZE (D_SIZE),
    .LOW_WIDTH (LOW_WIDTH),
    .RANGE_WIDTH (RANGE_WIDTH)
    ) s3_cdf (
      .u (u),
      .in_d (d),
      .in_s (in_s),
      .in_low (in_low),
      .in_range (in_range),
      .COMP_mux_1 (COMP_mux_1),
      // Outputs
      .out_s (s_cdf),
      .out_low (low_cdf),
      .out_bit_1 (out_bit_1_cdf),
      .out_bit_2 (out_bit_2_cdf),
      .flag_bitstream (flag_cdf)
    );

    s3_bool #(
      .D_SIZE (D_SIZE),
      .LOW_WIDTH (LOW_WIDTH),
      .RANGE_WIDTH (RANGE_WIDTH)
      ) s3_bool (
        .in_d (d),
        .in_s (in_s),
        .in_low (in_low),
        .symbol (symbol),
        .pre_low (pre_low),
        .in_range (in_range),
        // Outputs
        .out_s (s_bool),
        .out_low (low_bool),
        .out_bit_1 (bool_out_bit_1),
        .out_bit_2 (bool_out_bit_2),
        .flag_bitstream (flag_bit_bool)
    );

  // ------------------------------------------------------
  assign out_low =  (bool_flag) ? low_bool :
                    low_cdf;
  assign out_s =  (bool_flag) ? s_bool :
                  s_cdf;
  assign flag_bitstream = (bool_flag) ? flag_bit_bool :
                          flag_cdf;
  assign out_bit_1 =  (bool_flag) ? bool_out_bit_1 :
                      out_bit_1_cdf;
  assign out_bit_2 =  (bool_flag) ? bool_out_bit_2 :
                      out_bit_2_cdf;
  // Assigned Outputs
  assign out_range = range_ready;
endmodule

module s3_cdf #(
  parameter D_SIZE = 5,
  parameter LOW_WIDTH = 24,
  parameter RANGE_WIDTH = 16
  )(
    input COMP_mux_1,
    input [RANGE_WIDTH:0] u,
    input [(LOW_WIDTH-1):0] in_low,
    input [(D_SIZE-1):0] in_d, in_s,
    input [(RANGE_WIDTH-1):0] in_range,
    // Outputs
    output wire [1:0] flag_bitstream,
    output wire [(D_SIZE-1):0] out_s,
    output wire [(LOW_WIDTH-1):0] out_low,
    output wire [(RANGE_WIDTH-1):0] out_bit_1, out_bit_2
  );
  wire [(LOW_WIDTH-1):0] low_1, low_raw;
  assign low_1 = in_low + (in_range - u[(RANGE_WIDTH-1):0]);

  assign low_raw =  (COMP_mux_1 == 1'b1) ? low_1 :
                    in_low;
  s3_renormalization # (
    .D_SIZE (D_SIZE),
    .LOW_WIDTH (LOW_WIDTH),
    .RANGE_WIDTH (RANGE_WIDTH)
    ) s3_cdf_norm (
      .d (in_d),
      .in_s (in_s),
      .low_raw (low_raw),
      // Outputs
      .out_s (out_s),
      .out_low (out_low),
      .out_bit_1 (out_bit_1),
      .out_bit_2 (out_bit_2),
      .flag_bitstream (flag_bitstream)
    );
endmodule

module s3_bool #(
  parameter D_SIZE = 5,
  parameter LOW_WIDTH = 24,
  parameter RANGE_WIDTH = 16
  )(
    input symbol,
    input [(LOW_WIDTH-1):0] in_low,
    input [(D_SIZE-1):0] in_d, in_s,
    input [(RANGE_WIDTH-1):0] in_range, pre_low,
    // Outputs
    output wire [1:0] flag_bitstream,
    output wire [(D_SIZE-1):0] out_s,
    output wire [(LOW_WIDTH-1):0] out_low,
    output wire [(RANGE_WIDTH-1):0] out_bit_1, out_bit_2
  );
  wire [(LOW_WIDTH-1):0] low_1, low_raw;
  /* Pre_low is a variable calculated within the Boolean block in Stage 2.
    Its creation was specifically done to reduce the stress generated by the
  parallelized Boolean blocks in Stage 3.
    Pre_low = in_range - v_bool
  */
  assign low_1 = in_low + pre_low;

  assign low_raw =  (symbol == 1'b1) ? low_1 :
                    in_low;
  s3_renormalization #(
    .D_SIZE (D_SIZE),
    .LOW_WIDTH (LOW_WIDTH),
    .RANGE_WIDTH (RANGE_WIDTH)
    ) s3_bool_norm (
      .d (in_d),
      .in_s (in_s),
      .low_raw (low_raw),
      // Outputs
      .out_s (out_s),
      .out_low (out_low),
      .out_bit_1 (out_bit_1),
      .out_bit_2 (out_bit_2),
      .flag_bitstream (flag_bitstream)
    );
endmodule

module s3_renormalization #(
  parameter LOW_WIDTH = 24,
  parameter RANGE_WIDTH = 16,
  parameter D_SIZE = 5
  )(
    input [(LOW_WIDTH-1):0] low_raw,
    input [(D_SIZE-1):0] d, in_s,
    // Outputs
    output wire [1:0] flag_bitstream,
    output wire [(D_SIZE-1):0] out_s,
    output wire [(LOW_WIDTH-1):0] out_low,
    output wire [(RANGE_WIDTH-1):0] out_bit_1, out_bit_2
  );
  wire [(LOW_WIDTH-1):0] low_s0, low_s8, m_s8, m_s0;
  wire [(D_SIZE-1):0] c_norm_s0, c_norm_s8, s_s0, s_s8;
  wire [(D_SIZE-1):0] s_comp;
  wire [(D_SIZE-1):0] c_bit_s0, c_bit_s8;

  assign s_comp = in_s + d;
  // ----------------------
  assign c_norm_s0 = in_s + 5'd7;
  assign m_s0 = (24'd1 << c_norm_s0) - 24'd1;

  // s_s0 adapted from: s0 = (in_s + 16) + d - 24
  assign s_s0 = in_s + d - 5'd8;
  assign low_s0 = low_raw & m_s0;
  // -----------------------
  assign c_norm_s8 = in_s - 5'd1;
  // m_s8 adapted from: m_s8 = m_s0 >> 8
  assign m_s8 = (24'd1 << c_norm_s8) - 24'd1;

  // s_s8 adapted from: s8 = (in_s + 8) + d - 24
  assign s_s8 = in_s + d - 5'd16;
  assign low_s8 = low_raw & m_s8;

  // pre-bitstream generation
  assign c_bit_s0 = in_s + 5'd7;
  assign c_bit_s8 = in_s - 5'd1;
  // =========================================================================
  // Outputs

  assign out_low =  ((s_comp >= 9) && (s_comp < 17)) ? low_s0 << d :
                    (s_comp >= 17) ? low_s8 << d :
                    low_raw << d;

  assign out_s =  ((s_comp >= 9) && (s_comp < 17)) ? s_s0 :
                  (s_comp >= 17) ? s_s8 :
                  s_comp;
  /*
    out_bit_1 and out_bit_2 are the pre-bitstreams generated by Stage 3.
    They are send to Stage 4 (carry propagation) for a reduction from a 9-bit to
  an 8-bit array.
  */
  assign out_bit_1 =  (s_comp >= 9) ? low_raw >> c_bit_s0 :
                      16'd0;
  assign out_bit_2 =  (s_comp >= 17) ? low_s0 >> c_bit_s8 :
                      16'd0;
  /*
  flag_bitstream represents how many pre-bitstreams are being in a given round
      01 (1): generating only out_bit_1
      10 (2): generating out_bit_1 and out_bit_2
  */

  assign flag_bitstream = ((s_comp >= 9) && (s_comp < 17)) ? 2'd1 :
                          (s_comp >= 17) ? 2'd2 :
                          2'd0;
endmodule
